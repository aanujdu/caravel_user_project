magic
tech sky130A
magscale 1 2
timestamp 1647724974
<< obsli1 >>
rect 1104 2159 138644 139281
<< obsm1 >>
rect 14 1244 139734 139312
<< metal2 >>
rect 662 141167 718 141967
rect 1950 141167 2006 141967
rect 3882 141167 3938 141967
rect 5170 141167 5226 141967
rect 6458 141167 6514 141967
rect 7746 141167 7802 141967
rect 9034 141167 9090 141967
rect 10322 141167 10378 141967
rect 11610 141167 11666 141967
rect 12898 141167 12954 141967
rect 14186 141167 14242 141967
rect 15474 141167 15530 141967
rect 16762 141167 16818 141967
rect 18694 141167 18750 141967
rect 19982 141167 20038 141967
rect 21270 141167 21326 141967
rect 22558 141167 22614 141967
rect 23846 141167 23902 141967
rect 25134 141167 25190 141967
rect 26422 141167 26478 141967
rect 27710 141167 27766 141967
rect 28998 141167 29054 141967
rect 30286 141167 30342 141967
rect 31574 141167 31630 141967
rect 33506 141167 33562 141967
rect 34794 141167 34850 141967
rect 36082 141167 36138 141967
rect 37370 141167 37426 141967
rect 38658 141167 38714 141967
rect 39946 141167 40002 141967
rect 41234 141167 41290 141967
rect 42522 141167 42578 141967
rect 43810 141167 43866 141967
rect 45098 141167 45154 141967
rect 46386 141167 46442 141967
rect 47674 141167 47730 141967
rect 49606 141167 49662 141967
rect 50894 141167 50950 141967
rect 52182 141167 52238 141967
rect 53470 141167 53526 141967
rect 54758 141167 54814 141967
rect 56046 141167 56102 141967
rect 57334 141167 57390 141967
rect 58622 141167 58678 141967
rect 59910 141167 59966 141967
rect 61198 141167 61254 141967
rect 62486 141167 62542 141967
rect 64418 141167 64474 141967
rect 65706 141167 65762 141967
rect 66994 141167 67050 141967
rect 68282 141167 68338 141967
rect 69570 141167 69626 141967
rect 70858 141167 70914 141967
rect 72146 141167 72202 141967
rect 73434 141167 73490 141967
rect 74722 141167 74778 141967
rect 76010 141167 76066 141967
rect 77298 141167 77354 141967
rect 78586 141167 78642 141967
rect 80518 141167 80574 141967
rect 81806 141167 81862 141967
rect 83094 141167 83150 141967
rect 84382 141167 84438 141967
rect 85670 141167 85726 141967
rect 86958 141167 87014 141967
rect 88246 141167 88302 141967
rect 89534 141167 89590 141967
rect 90822 141167 90878 141967
rect 92110 141167 92166 141967
rect 93398 141167 93454 141967
rect 95330 141167 95386 141967
rect 96618 141167 96674 141967
rect 97906 141167 97962 141967
rect 99194 141167 99250 141967
rect 100482 141167 100538 141967
rect 101770 141167 101826 141967
rect 103058 141167 103114 141967
rect 104346 141167 104402 141967
rect 105634 141167 105690 141967
rect 106922 141167 106978 141967
rect 108210 141167 108266 141967
rect 110142 141167 110198 141967
rect 111430 141167 111486 141967
rect 112718 141167 112774 141967
rect 114006 141167 114062 141967
rect 115294 141167 115350 141967
rect 116582 141167 116638 141967
rect 117870 141167 117926 141967
rect 119158 141167 119214 141967
rect 120446 141167 120502 141967
rect 121734 141167 121790 141967
rect 123022 141167 123078 141967
rect 124310 141167 124366 141967
rect 126242 141167 126298 141967
rect 127530 141167 127586 141967
rect 128818 141167 128874 141967
rect 130106 141167 130162 141967
rect 131394 141167 131450 141967
rect 132682 141167 132738 141967
rect 133970 141167 134026 141967
rect 135258 141167 135314 141967
rect 136546 141167 136602 141967
rect 137834 141167 137890 141967
rect 139122 141167 139178 141967
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 30930 0 30986 800
rect 32218 0 32274 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 45098 0 45154 800
rect 47030 0 47086 800
rect 48318 0 48374 800
rect 49606 0 49662 800
rect 50894 0 50950 800
rect 52182 0 52238 800
rect 53470 0 53526 800
rect 54758 0 54814 800
rect 56046 0 56102 800
rect 57334 0 57390 800
rect 58622 0 58678 800
rect 59910 0 59966 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 64418 0 64474 800
rect 65706 0 65762 800
rect 66994 0 67050 800
rect 68282 0 68338 800
rect 69570 0 69626 800
rect 70858 0 70914 800
rect 72146 0 72202 800
rect 73434 0 73490 800
rect 74722 0 74778 800
rect 76654 0 76710 800
rect 77942 0 77998 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 84382 0 84438 800
rect 85670 0 85726 800
rect 86958 0 87014 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 90822 0 90878 800
rect 92754 0 92810 800
rect 94042 0 94098 800
rect 95330 0 95386 800
rect 96618 0 96674 800
rect 97906 0 97962 800
rect 99194 0 99250 800
rect 100482 0 100538 800
rect 101770 0 101826 800
rect 103058 0 103114 800
rect 104346 0 104402 800
rect 105634 0 105690 800
rect 107566 0 107622 800
rect 108854 0 108910 800
rect 110142 0 110198 800
rect 111430 0 111486 800
rect 112718 0 112774 800
rect 114006 0 114062 800
rect 115294 0 115350 800
rect 116582 0 116638 800
rect 117870 0 117926 800
rect 119158 0 119214 800
rect 120446 0 120502 800
rect 122378 0 122434 800
rect 123666 0 123722 800
rect 124954 0 125010 800
rect 126242 0 126298 800
rect 127530 0 127586 800
rect 128818 0 128874 800
rect 130106 0 130162 800
rect 131394 0 131450 800
rect 132682 0 132738 800
rect 133970 0 134026 800
rect 135258 0 135314 800
rect 136546 0 136602 800
rect 138478 0 138534 800
rect 139766 0 139822 800
<< obsm2 >>
rect 20 141111 606 141545
rect 774 141111 1894 141545
rect 2062 141111 3826 141545
rect 3994 141111 5114 141545
rect 5282 141111 6402 141545
rect 6570 141111 7690 141545
rect 7858 141111 8978 141545
rect 9146 141111 10266 141545
rect 10434 141111 11554 141545
rect 11722 141111 12842 141545
rect 13010 141111 14130 141545
rect 14298 141111 15418 141545
rect 15586 141111 16706 141545
rect 16874 141111 18638 141545
rect 18806 141111 19926 141545
rect 20094 141111 21214 141545
rect 21382 141111 22502 141545
rect 22670 141111 23790 141545
rect 23958 141111 25078 141545
rect 25246 141111 26366 141545
rect 26534 141111 27654 141545
rect 27822 141111 28942 141545
rect 29110 141111 30230 141545
rect 30398 141111 31518 141545
rect 31686 141111 33450 141545
rect 33618 141111 34738 141545
rect 34906 141111 36026 141545
rect 36194 141111 37314 141545
rect 37482 141111 38602 141545
rect 38770 141111 39890 141545
rect 40058 141111 41178 141545
rect 41346 141111 42466 141545
rect 42634 141111 43754 141545
rect 43922 141111 45042 141545
rect 45210 141111 46330 141545
rect 46498 141111 47618 141545
rect 47786 141111 49550 141545
rect 49718 141111 50838 141545
rect 51006 141111 52126 141545
rect 52294 141111 53414 141545
rect 53582 141111 54702 141545
rect 54870 141111 55990 141545
rect 56158 141111 57278 141545
rect 57446 141111 58566 141545
rect 58734 141111 59854 141545
rect 60022 141111 61142 141545
rect 61310 141111 62430 141545
rect 62598 141111 64362 141545
rect 64530 141111 65650 141545
rect 65818 141111 66938 141545
rect 67106 141111 68226 141545
rect 68394 141111 69514 141545
rect 69682 141111 70802 141545
rect 70970 141111 72090 141545
rect 72258 141111 73378 141545
rect 73546 141111 74666 141545
rect 74834 141111 75954 141545
rect 76122 141111 77242 141545
rect 77410 141111 78530 141545
rect 78698 141111 80462 141545
rect 80630 141111 81750 141545
rect 81918 141111 83038 141545
rect 83206 141111 84326 141545
rect 84494 141111 85614 141545
rect 85782 141111 86902 141545
rect 87070 141111 88190 141545
rect 88358 141111 89478 141545
rect 89646 141111 90766 141545
rect 90934 141111 92054 141545
rect 92222 141111 93342 141545
rect 93510 141111 95274 141545
rect 95442 141111 96562 141545
rect 96730 141111 97850 141545
rect 98018 141111 99138 141545
rect 99306 141111 100426 141545
rect 100594 141111 101714 141545
rect 101882 141111 103002 141545
rect 103170 141111 104290 141545
rect 104458 141111 105578 141545
rect 105746 141111 106866 141545
rect 107034 141111 108154 141545
rect 108322 141111 110086 141545
rect 110254 141111 111374 141545
rect 111542 141111 112662 141545
rect 112830 141111 113950 141545
rect 114118 141111 115238 141545
rect 115406 141111 116526 141545
rect 116694 141111 117814 141545
rect 117982 141111 119102 141545
rect 119270 141111 120390 141545
rect 120558 141111 121678 141545
rect 121846 141111 122966 141545
rect 123134 141111 124254 141545
rect 124422 141111 126186 141545
rect 126354 141111 127474 141545
rect 127642 141111 128762 141545
rect 128930 141111 130050 141545
rect 130218 141111 131338 141545
rect 131506 141111 132626 141545
rect 132794 141111 133914 141545
rect 134082 141111 135202 141545
rect 135370 141111 136490 141545
rect 136658 141111 137778 141545
rect 137946 141111 139066 141545
rect 139234 141111 139808 141545
rect 20 856 139808 141111
rect 130 734 1250 856
rect 1418 734 2538 856
rect 2706 734 3826 856
rect 3994 734 5114 856
rect 5282 734 6402 856
rect 6570 734 7690 856
rect 7858 734 8978 856
rect 9146 734 10266 856
rect 10434 734 11554 856
rect 11722 734 12842 856
rect 13010 734 14130 856
rect 14298 734 16062 856
rect 16230 734 17350 856
rect 17518 734 18638 856
rect 18806 734 19926 856
rect 20094 734 21214 856
rect 21382 734 22502 856
rect 22670 734 23790 856
rect 23958 734 25078 856
rect 25246 734 26366 856
rect 26534 734 27654 856
rect 27822 734 28942 856
rect 29110 734 30874 856
rect 31042 734 32162 856
rect 32330 734 33450 856
rect 33618 734 34738 856
rect 34906 734 36026 856
rect 36194 734 37314 856
rect 37482 734 38602 856
rect 38770 734 39890 856
rect 40058 734 41178 856
rect 41346 734 42466 856
rect 42634 734 43754 856
rect 43922 734 45042 856
rect 45210 734 46974 856
rect 47142 734 48262 856
rect 48430 734 49550 856
rect 49718 734 50838 856
rect 51006 734 52126 856
rect 52294 734 53414 856
rect 53582 734 54702 856
rect 54870 734 55990 856
rect 56158 734 57278 856
rect 57446 734 58566 856
rect 58734 734 59854 856
rect 60022 734 61786 856
rect 61954 734 63074 856
rect 63242 734 64362 856
rect 64530 734 65650 856
rect 65818 734 66938 856
rect 67106 734 68226 856
rect 68394 734 69514 856
rect 69682 734 70802 856
rect 70970 734 72090 856
rect 72258 734 73378 856
rect 73546 734 74666 856
rect 74834 734 76598 856
rect 76766 734 77886 856
rect 78054 734 79174 856
rect 79342 734 80462 856
rect 80630 734 81750 856
rect 81918 734 83038 856
rect 83206 734 84326 856
rect 84494 734 85614 856
rect 85782 734 86902 856
rect 87070 734 88190 856
rect 88358 734 89478 856
rect 89646 734 90766 856
rect 90934 734 92698 856
rect 92866 734 93986 856
rect 94154 734 95274 856
rect 95442 734 96562 856
rect 96730 734 97850 856
rect 98018 734 99138 856
rect 99306 734 100426 856
rect 100594 734 101714 856
rect 101882 734 103002 856
rect 103170 734 104290 856
rect 104458 734 105578 856
rect 105746 734 107510 856
rect 107678 734 108798 856
rect 108966 734 110086 856
rect 110254 734 111374 856
rect 111542 734 112662 856
rect 112830 734 113950 856
rect 114118 734 115238 856
rect 115406 734 116526 856
rect 116694 734 117814 856
rect 117982 734 119102 856
rect 119270 734 120390 856
rect 120558 734 122322 856
rect 122490 734 123610 856
rect 123778 734 124898 856
rect 125066 734 126186 856
rect 126354 734 127474 856
rect 127642 734 128762 856
rect 128930 734 130050 856
rect 130218 734 131338 856
rect 131506 734 132626 856
rect 132794 734 133914 856
rect 134082 734 135202 856
rect 135370 734 136490 856
rect 136658 734 138422 856
rect 138590 734 139710 856
<< metal3 >>
rect 0 141448 800 141568
rect 139023 140768 139823 140888
rect 0 140088 800 140208
rect 139023 139408 139823 139528
rect 0 138728 800 138848
rect 139023 138048 139823 138168
rect 0 137368 800 137488
rect 139023 136688 139823 136808
rect 0 136008 800 136128
rect 139023 135328 139823 135448
rect 0 134648 800 134768
rect 139023 133968 139823 134088
rect 0 133288 800 133408
rect 139023 132608 139823 132728
rect 0 131928 800 132048
rect 139023 131248 139823 131368
rect 0 130568 800 130688
rect 139023 129888 139823 130008
rect 0 129208 800 129328
rect 139023 128528 139823 128648
rect 0 127168 800 127288
rect 139023 127168 139823 127288
rect 0 125808 800 125928
rect 139023 125128 139823 125248
rect 0 124448 800 124568
rect 139023 123768 139823 123888
rect 0 123088 800 123208
rect 139023 122408 139823 122528
rect 0 121728 800 121848
rect 139023 121048 139823 121168
rect 0 120368 800 120488
rect 139023 119688 139823 119808
rect 0 119008 800 119128
rect 139023 118328 139823 118448
rect 0 117648 800 117768
rect 139023 116968 139823 117088
rect 0 116288 800 116408
rect 139023 115608 139823 115728
rect 0 114928 800 115048
rect 139023 114248 139823 114368
rect 0 113568 800 113688
rect 139023 112888 139823 113008
rect 0 111528 800 111648
rect 139023 111528 139823 111648
rect 0 110168 800 110288
rect 139023 110168 139823 110288
rect 0 108808 800 108928
rect 139023 108128 139823 108248
rect 0 107448 800 107568
rect 139023 106768 139823 106888
rect 0 106088 800 106208
rect 139023 105408 139823 105528
rect 0 104728 800 104848
rect 139023 104048 139823 104168
rect 0 103368 800 103488
rect 139023 102688 139823 102808
rect 0 102008 800 102128
rect 139023 101328 139823 101448
rect 0 100648 800 100768
rect 139023 99968 139823 100088
rect 0 99288 800 99408
rect 139023 98608 139823 98728
rect 0 97928 800 98048
rect 139023 97248 139823 97368
rect 0 95888 800 96008
rect 139023 95888 139823 96008
rect 0 94528 800 94648
rect 139023 94528 139823 94648
rect 0 93168 800 93288
rect 139023 92488 139823 92608
rect 0 91808 800 91928
rect 139023 91128 139823 91248
rect 0 90448 800 90568
rect 139023 89768 139823 89888
rect 0 89088 800 89208
rect 139023 88408 139823 88528
rect 0 87728 800 87848
rect 139023 87048 139823 87168
rect 0 86368 800 86488
rect 139023 85688 139823 85808
rect 0 85008 800 85128
rect 139023 84328 139823 84448
rect 0 83648 800 83768
rect 139023 82968 139823 83088
rect 0 82288 800 82408
rect 139023 81608 139823 81728
rect 0 80928 800 81048
rect 139023 80248 139823 80368
rect 0 78888 800 79008
rect 139023 78888 139823 79008
rect 0 77528 800 77648
rect 139023 76848 139823 76968
rect 0 76168 800 76288
rect 139023 75488 139823 75608
rect 0 74808 800 74928
rect 139023 74128 139823 74248
rect 0 73448 800 73568
rect 139023 72768 139823 72888
rect 0 72088 800 72208
rect 139023 71408 139823 71528
rect 0 70728 800 70848
rect 139023 70048 139823 70168
rect 0 69368 800 69488
rect 139023 68688 139823 68808
rect 0 68008 800 68128
rect 139023 67328 139823 67448
rect 0 66648 800 66768
rect 139023 65968 139823 66088
rect 0 65288 800 65408
rect 139023 64608 139823 64728
rect 0 63248 800 63368
rect 139023 63248 139823 63368
rect 0 61888 800 62008
rect 139023 61888 139823 62008
rect 0 60528 800 60648
rect 139023 59848 139823 59968
rect 0 59168 800 59288
rect 139023 58488 139823 58608
rect 0 57808 800 57928
rect 139023 57128 139823 57248
rect 0 56448 800 56568
rect 139023 55768 139823 55888
rect 0 55088 800 55208
rect 139023 54408 139823 54528
rect 0 53728 800 53848
rect 139023 53048 139823 53168
rect 0 52368 800 52488
rect 139023 51688 139823 51808
rect 0 51008 800 51128
rect 139023 50328 139823 50448
rect 0 49648 800 49768
rect 139023 48968 139823 49088
rect 0 47608 800 47728
rect 139023 47608 139823 47728
rect 0 46248 800 46368
rect 139023 46248 139823 46368
rect 0 44888 800 45008
rect 139023 44208 139823 44328
rect 0 43528 800 43648
rect 139023 42848 139823 42968
rect 0 42168 800 42288
rect 139023 41488 139823 41608
rect 0 40808 800 40928
rect 139023 40128 139823 40248
rect 0 39448 800 39568
rect 139023 38768 139823 38888
rect 0 38088 800 38208
rect 139023 37408 139823 37528
rect 0 36728 800 36848
rect 139023 36048 139823 36168
rect 0 35368 800 35488
rect 139023 34688 139823 34808
rect 0 34008 800 34128
rect 139023 33328 139823 33448
rect 0 32648 800 32768
rect 139023 31968 139823 32088
rect 0 30608 800 30728
rect 139023 30608 139823 30728
rect 0 29248 800 29368
rect 139023 29248 139823 29368
rect 0 27888 800 28008
rect 139023 27208 139823 27328
rect 0 26528 800 26648
rect 139023 25848 139823 25968
rect 0 25168 800 25288
rect 139023 24488 139823 24608
rect 0 23808 800 23928
rect 139023 23128 139823 23248
rect 0 22448 800 22568
rect 139023 21768 139823 21888
rect 0 21088 800 21208
rect 139023 20408 139823 20528
rect 0 19728 800 19848
rect 139023 19048 139823 19168
rect 0 18368 800 18488
rect 139023 17688 139823 17808
rect 0 17008 800 17128
rect 139023 16328 139823 16448
rect 0 14968 800 15088
rect 139023 14968 139823 15088
rect 0 13608 800 13728
rect 139023 13608 139823 13728
rect 0 12248 800 12368
rect 139023 11568 139823 11688
rect 0 10888 800 11008
rect 139023 10208 139823 10328
rect 0 9528 800 9648
rect 139023 8848 139823 8968
rect 0 8168 800 8288
rect 139023 7488 139823 7608
rect 0 6808 800 6928
rect 139023 6128 139823 6248
rect 0 5448 800 5568
rect 139023 4768 139823 4888
rect 0 4088 800 4208
rect 139023 3408 139823 3528
rect 0 2728 800 2848
rect 139023 2048 139823 2168
rect 0 1368 800 1488
rect 139023 688 139823 808
<< obsm3 >>
rect 880 141368 139023 141541
rect 565 140968 139023 141368
rect 565 140688 138943 140968
rect 565 140288 139023 140688
rect 880 140008 139023 140288
rect 565 139608 139023 140008
rect 565 139328 138943 139608
rect 565 138928 139023 139328
rect 880 138648 139023 138928
rect 565 138248 139023 138648
rect 565 137968 138943 138248
rect 565 137568 139023 137968
rect 880 137288 139023 137568
rect 565 136888 139023 137288
rect 565 136608 138943 136888
rect 565 136208 139023 136608
rect 880 135928 139023 136208
rect 565 135528 139023 135928
rect 565 135248 138943 135528
rect 565 134848 139023 135248
rect 880 134568 139023 134848
rect 565 134168 139023 134568
rect 565 133888 138943 134168
rect 565 133488 139023 133888
rect 880 133208 139023 133488
rect 565 132808 139023 133208
rect 565 132528 138943 132808
rect 565 132128 139023 132528
rect 880 131848 139023 132128
rect 565 131448 139023 131848
rect 565 131168 138943 131448
rect 565 130768 139023 131168
rect 880 130488 139023 130768
rect 565 130088 139023 130488
rect 565 129808 138943 130088
rect 565 129408 139023 129808
rect 880 129128 139023 129408
rect 565 128728 139023 129128
rect 565 128448 138943 128728
rect 565 127368 139023 128448
rect 880 127088 138943 127368
rect 565 126008 139023 127088
rect 880 125728 139023 126008
rect 565 125328 139023 125728
rect 565 125048 138943 125328
rect 565 124648 139023 125048
rect 880 124368 139023 124648
rect 565 123968 139023 124368
rect 565 123688 138943 123968
rect 565 123288 139023 123688
rect 880 123008 139023 123288
rect 565 122608 139023 123008
rect 565 122328 138943 122608
rect 565 121928 139023 122328
rect 880 121648 139023 121928
rect 565 121248 139023 121648
rect 565 120968 138943 121248
rect 565 120568 139023 120968
rect 880 120288 139023 120568
rect 565 119888 139023 120288
rect 565 119608 138943 119888
rect 565 119208 139023 119608
rect 880 118928 139023 119208
rect 565 118528 139023 118928
rect 565 118248 138943 118528
rect 565 117848 139023 118248
rect 880 117568 139023 117848
rect 565 117168 139023 117568
rect 565 116888 138943 117168
rect 565 116488 139023 116888
rect 880 116208 139023 116488
rect 565 115808 139023 116208
rect 565 115528 138943 115808
rect 565 115128 139023 115528
rect 880 114848 139023 115128
rect 565 114448 139023 114848
rect 565 114168 138943 114448
rect 565 113768 139023 114168
rect 880 113488 139023 113768
rect 565 113088 139023 113488
rect 565 112808 138943 113088
rect 565 111728 139023 112808
rect 880 111448 138943 111728
rect 565 110368 139023 111448
rect 880 110088 138943 110368
rect 565 109008 139023 110088
rect 880 108728 139023 109008
rect 565 108328 139023 108728
rect 565 108048 138943 108328
rect 565 107648 139023 108048
rect 880 107368 139023 107648
rect 565 106968 139023 107368
rect 565 106688 138943 106968
rect 565 106288 139023 106688
rect 880 106008 139023 106288
rect 565 105608 139023 106008
rect 565 105328 138943 105608
rect 565 104928 139023 105328
rect 880 104648 139023 104928
rect 565 104248 139023 104648
rect 565 103968 138943 104248
rect 565 103568 139023 103968
rect 880 103288 139023 103568
rect 565 102888 139023 103288
rect 565 102608 138943 102888
rect 565 102208 139023 102608
rect 880 101928 139023 102208
rect 565 101528 139023 101928
rect 565 101248 138943 101528
rect 565 100848 139023 101248
rect 880 100568 139023 100848
rect 565 100168 139023 100568
rect 565 99888 138943 100168
rect 565 99488 139023 99888
rect 880 99208 139023 99488
rect 565 98808 139023 99208
rect 565 98528 138943 98808
rect 565 98128 139023 98528
rect 880 97848 139023 98128
rect 565 97448 139023 97848
rect 565 97168 138943 97448
rect 565 96088 139023 97168
rect 880 95808 138943 96088
rect 565 94728 139023 95808
rect 880 94448 138943 94728
rect 565 93368 139023 94448
rect 880 93088 139023 93368
rect 565 92688 139023 93088
rect 565 92408 138943 92688
rect 565 92008 139023 92408
rect 880 91728 139023 92008
rect 565 91328 139023 91728
rect 565 91048 138943 91328
rect 565 90648 139023 91048
rect 880 90368 139023 90648
rect 565 89968 139023 90368
rect 565 89688 138943 89968
rect 565 89288 139023 89688
rect 880 89008 139023 89288
rect 565 88608 139023 89008
rect 565 88328 138943 88608
rect 565 87928 139023 88328
rect 880 87648 139023 87928
rect 565 87248 139023 87648
rect 565 86968 138943 87248
rect 565 86568 139023 86968
rect 880 86288 139023 86568
rect 565 85888 139023 86288
rect 565 85608 138943 85888
rect 565 85208 139023 85608
rect 880 84928 139023 85208
rect 565 84528 139023 84928
rect 565 84248 138943 84528
rect 565 83848 139023 84248
rect 880 83568 139023 83848
rect 565 83168 139023 83568
rect 565 82888 138943 83168
rect 565 82488 139023 82888
rect 880 82208 139023 82488
rect 565 81808 139023 82208
rect 565 81528 138943 81808
rect 565 81128 139023 81528
rect 880 80848 139023 81128
rect 565 80448 139023 80848
rect 565 80168 138943 80448
rect 565 79088 139023 80168
rect 880 78808 138943 79088
rect 565 77728 139023 78808
rect 880 77448 139023 77728
rect 565 77048 139023 77448
rect 565 76768 138943 77048
rect 565 76368 139023 76768
rect 880 76088 139023 76368
rect 565 75688 139023 76088
rect 565 75408 138943 75688
rect 565 75008 139023 75408
rect 880 74728 139023 75008
rect 565 74328 139023 74728
rect 565 74048 138943 74328
rect 565 73648 139023 74048
rect 880 73368 139023 73648
rect 565 72968 139023 73368
rect 565 72688 138943 72968
rect 565 72288 139023 72688
rect 880 72008 139023 72288
rect 565 71608 139023 72008
rect 565 71328 138943 71608
rect 565 70928 139023 71328
rect 880 70648 139023 70928
rect 565 70248 139023 70648
rect 565 69968 138943 70248
rect 565 69568 139023 69968
rect 880 69288 139023 69568
rect 565 68888 139023 69288
rect 565 68608 138943 68888
rect 565 68208 139023 68608
rect 880 67928 139023 68208
rect 565 67528 139023 67928
rect 565 67248 138943 67528
rect 565 66848 139023 67248
rect 880 66568 139023 66848
rect 565 66168 139023 66568
rect 565 65888 138943 66168
rect 565 65488 139023 65888
rect 880 65208 139023 65488
rect 565 64808 139023 65208
rect 565 64528 138943 64808
rect 565 63448 139023 64528
rect 880 63168 138943 63448
rect 565 62088 139023 63168
rect 880 61808 138943 62088
rect 565 60728 139023 61808
rect 880 60448 139023 60728
rect 565 60048 139023 60448
rect 565 59768 138943 60048
rect 565 59368 139023 59768
rect 880 59088 139023 59368
rect 565 58688 139023 59088
rect 565 58408 138943 58688
rect 565 58008 139023 58408
rect 880 57728 139023 58008
rect 565 57328 139023 57728
rect 565 57048 138943 57328
rect 565 56648 139023 57048
rect 880 56368 139023 56648
rect 565 55968 139023 56368
rect 565 55688 138943 55968
rect 565 55288 139023 55688
rect 880 55008 139023 55288
rect 565 54608 139023 55008
rect 565 54328 138943 54608
rect 565 53928 139023 54328
rect 880 53648 139023 53928
rect 565 53248 139023 53648
rect 565 52968 138943 53248
rect 565 52568 139023 52968
rect 880 52288 139023 52568
rect 565 51888 139023 52288
rect 565 51608 138943 51888
rect 565 51208 139023 51608
rect 880 50928 139023 51208
rect 565 50528 139023 50928
rect 565 50248 138943 50528
rect 565 49848 139023 50248
rect 880 49568 139023 49848
rect 565 49168 139023 49568
rect 565 48888 138943 49168
rect 565 47808 139023 48888
rect 880 47528 138943 47808
rect 565 46448 139023 47528
rect 880 46168 138943 46448
rect 565 45088 139023 46168
rect 880 44808 139023 45088
rect 565 44408 139023 44808
rect 565 44128 138943 44408
rect 565 43728 139023 44128
rect 880 43448 139023 43728
rect 565 43048 139023 43448
rect 565 42768 138943 43048
rect 565 42368 139023 42768
rect 880 42088 139023 42368
rect 565 41688 139023 42088
rect 565 41408 138943 41688
rect 565 41008 139023 41408
rect 880 40728 139023 41008
rect 565 40328 139023 40728
rect 565 40048 138943 40328
rect 565 39648 139023 40048
rect 880 39368 139023 39648
rect 565 38968 139023 39368
rect 565 38688 138943 38968
rect 565 38288 139023 38688
rect 880 38008 139023 38288
rect 565 37608 139023 38008
rect 565 37328 138943 37608
rect 565 36928 139023 37328
rect 880 36648 139023 36928
rect 565 36248 139023 36648
rect 565 35968 138943 36248
rect 565 35568 139023 35968
rect 880 35288 139023 35568
rect 565 34888 139023 35288
rect 565 34608 138943 34888
rect 565 34208 139023 34608
rect 880 33928 139023 34208
rect 565 33528 139023 33928
rect 565 33248 138943 33528
rect 565 32848 139023 33248
rect 880 32568 139023 32848
rect 565 32168 139023 32568
rect 565 31888 138943 32168
rect 565 30808 139023 31888
rect 880 30528 138943 30808
rect 565 29448 139023 30528
rect 880 29168 138943 29448
rect 565 28088 139023 29168
rect 880 27808 139023 28088
rect 565 27408 139023 27808
rect 565 27128 138943 27408
rect 565 26728 139023 27128
rect 880 26448 139023 26728
rect 565 26048 139023 26448
rect 565 25768 138943 26048
rect 565 25368 139023 25768
rect 880 25088 139023 25368
rect 565 24688 139023 25088
rect 565 24408 138943 24688
rect 565 24008 139023 24408
rect 880 23728 139023 24008
rect 565 23328 139023 23728
rect 565 23048 138943 23328
rect 565 22648 139023 23048
rect 880 22368 139023 22648
rect 565 21968 139023 22368
rect 565 21688 138943 21968
rect 565 21288 139023 21688
rect 880 21008 139023 21288
rect 565 20608 139023 21008
rect 565 20328 138943 20608
rect 565 19928 139023 20328
rect 880 19648 139023 19928
rect 565 19248 139023 19648
rect 565 18968 138943 19248
rect 565 18568 139023 18968
rect 880 18288 139023 18568
rect 565 17888 139023 18288
rect 565 17608 138943 17888
rect 565 17208 139023 17608
rect 880 16928 139023 17208
rect 565 16528 139023 16928
rect 565 16248 138943 16528
rect 565 15168 139023 16248
rect 880 14888 138943 15168
rect 565 13808 139023 14888
rect 880 13528 138943 13808
rect 565 12448 139023 13528
rect 880 12168 139023 12448
rect 565 11768 139023 12168
rect 565 11488 138943 11768
rect 565 11088 139023 11488
rect 880 10808 139023 11088
rect 565 10408 139023 10808
rect 565 10128 138943 10408
rect 565 9728 139023 10128
rect 880 9448 139023 9728
rect 565 9048 139023 9448
rect 565 8768 138943 9048
rect 565 8368 139023 8768
rect 880 8088 139023 8368
rect 565 7688 139023 8088
rect 565 7408 138943 7688
rect 565 7008 139023 7408
rect 880 6728 139023 7008
rect 565 6328 139023 6728
rect 565 6048 138943 6328
rect 565 5648 139023 6048
rect 880 5368 139023 5648
rect 565 4968 139023 5368
rect 565 4688 138943 4968
rect 565 4288 139023 4688
rect 880 4008 139023 4288
rect 565 3608 139023 4008
rect 565 3328 138943 3608
rect 565 2928 139023 3328
rect 880 2648 139023 2928
rect 565 2248 139023 2648
rect 565 1968 138943 2248
rect 565 1568 139023 1968
rect 880 1288 139023 1568
rect 565 888 139023 1288
rect 565 718 138943 888
<< metal4 >>
rect 4208 2128 4528 139312
rect 19568 2128 19888 139312
rect 34928 2128 35248 139312
rect 50288 2128 50608 139312
rect 65648 2128 65968 139312
rect 81008 2128 81328 139312
rect 96368 2128 96688 139312
rect 111728 2128 112048 139312
rect 127088 2128 127408 139312
<< obsm4 >>
rect 1899 2048 4128 138141
rect 4608 2048 19488 138141
rect 19968 2048 34848 138141
rect 35328 2048 50208 138141
rect 50688 2048 65568 138141
rect 66048 2048 80928 138141
rect 81408 2048 96288 138141
rect 96768 2048 111648 138141
rect 112128 2048 127008 138141
rect 127488 2048 137573 138141
rect 1899 1395 137573 2048
<< obsm5 >>
rect 2508 37580 70540 56940
<< labels >>
rlabel metal4 s 19568 2128 19888 139312 6 VGND
port 1 nsew ground input
rlabel metal4 s 50288 2128 50608 139312 6 VGND
port 1 nsew ground input
rlabel metal4 s 81008 2128 81328 139312 6 VGND
port 1 nsew ground input
rlabel metal4 s 111728 2128 112048 139312 6 VGND
port 1 nsew ground input
rlabel metal4 s 4208 2128 4528 139312 6 VPWR
port 2 nsew power input
rlabel metal4 s 34928 2128 35248 139312 6 VPWR
port 2 nsew power input
rlabel metal4 s 65648 2128 65968 139312 6 VPWR
port 2 nsew power input
rlabel metal4 s 96368 2128 96688 139312 6 VPWR
port 2 nsew power input
rlabel metal4 s 127088 2128 127408 139312 6 VPWR
port 2 nsew power input
rlabel metal3 s 139023 136688 139823 136808 6 clk
port 3 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 eoi[0]
port 4 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 eoi[10]
port 5 nsew signal output
rlabel metal3 s 139023 8848 139823 8968 6 eoi[11]
port 6 nsew signal output
rlabel metal3 s 139023 88408 139823 88528 6 eoi[12]
port 7 nsew signal output
rlabel metal2 s 120446 141167 120502 141967 6 eoi[13]
port 8 nsew signal output
rlabel metal3 s 139023 74128 139823 74248 6 eoi[14]
port 9 nsew signal output
rlabel metal3 s 139023 23128 139823 23248 6 eoi[15]
port 10 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 eoi[16]
port 11 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 eoi[17]
port 12 nsew signal output
rlabel metal3 s 139023 17688 139823 17808 6 eoi[18]
port 13 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 eoi[19]
port 14 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 eoi[1]
port 15 nsew signal output
rlabel metal3 s 139023 64608 139823 64728 6 eoi[20]
port 16 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 eoi[21]
port 17 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 eoi[22]
port 18 nsew signal output
rlabel metal3 s 139023 25848 139823 25968 6 eoi[23]
port 19 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 eoi[24]
port 20 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 eoi[25]
port 21 nsew signal output
rlabel metal2 s 58622 141167 58678 141967 6 eoi[26]
port 22 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 eoi[27]
port 23 nsew signal output
rlabel metal3 s 139023 19048 139823 19168 6 eoi[28]
port 24 nsew signal output
rlabel metal3 s 139023 42848 139823 42968 6 eoi[29]
port 25 nsew signal output
rlabel metal3 s 139023 106768 139823 106888 6 eoi[2]
port 26 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 eoi[30]
port 27 nsew signal output
rlabel metal3 s 139023 72768 139823 72888 6 eoi[31]
port 28 nsew signal output
rlabel metal2 s 42522 141167 42578 141967 6 eoi[3]
port 29 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 eoi[4]
port 30 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 eoi[5]
port 31 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 eoi[6]
port 32 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 eoi[7]
port 33 nsew signal output
rlabel metal2 s 103058 141167 103114 141967 6 eoi[8]
port 34 nsew signal output
rlabel metal2 s 77298 141167 77354 141967 6 eoi[9]
port 35 nsew signal output
rlabel metal3 s 139023 55768 139823 55888 6 irq[0]
port 36 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 irq[10]
port 37 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 irq[11]
port 38 nsew signal input
rlabel metal2 s 85670 141167 85726 141967 6 irq[12]
port 39 nsew signal input
rlabel metal2 s 135258 141167 135314 141967 6 irq[13]
port 40 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 irq[14]
port 41 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 irq[15]
port 42 nsew signal input
rlabel metal2 s 139122 141167 139178 141967 6 irq[16]
port 43 nsew signal input
rlabel metal2 s 78586 141167 78642 141967 6 irq[17]
port 44 nsew signal input
rlabel metal2 s 105634 141167 105690 141967 6 irq[18]
port 45 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 irq[19]
port 46 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 irq[1]
port 47 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 irq[20]
port 48 nsew signal input
rlabel metal3 s 139023 85688 139823 85808 6 irq[21]
port 49 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 irq[22]
port 50 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 irq[23]
port 51 nsew signal input
rlabel metal3 s 139023 140768 139823 140888 6 irq[24]
port 52 nsew signal input
rlabel metal2 s 34794 141167 34850 141967 6 irq[25]
port 53 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 irq[26]
port 54 nsew signal input
rlabel metal2 s 70858 141167 70914 141967 6 irq[27]
port 55 nsew signal input
rlabel metal3 s 139023 133968 139823 134088 6 irq[28]
port 56 nsew signal input
rlabel metal3 s 139023 16328 139823 16448 6 irq[29]
port 57 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 irq[2]
port 58 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 irq[30]
port 59 nsew signal input
rlabel metal2 s 33506 141167 33562 141967 6 irq[31]
port 60 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 irq[3]
port 61 nsew signal input
rlabel metal2 s 27710 141167 27766 141967 6 irq[4]
port 62 nsew signal input
rlabel metal3 s 139023 125128 139823 125248 6 irq[5]
port 63 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 irq[6]
port 64 nsew signal input
rlabel metal2 s 3882 141167 3938 141967 6 irq[7]
port 65 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 irq[8]
port 66 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 irq[9]
port 67 nsew signal input
rlabel metal3 s 139023 3408 139823 3528 6 mem_addr[0]
port 68 nsew signal output
rlabel metal3 s 139023 67328 139823 67448 6 mem_addr[10]
port 69 nsew signal output
rlabel metal3 s 139023 121048 139823 121168 6 mem_addr[11]
port 70 nsew signal output
rlabel metal3 s 139023 14968 139823 15088 6 mem_addr[12]
port 71 nsew signal output
rlabel metal2 s 81806 141167 81862 141967 6 mem_addr[13]
port 72 nsew signal output
rlabel metal2 s 116582 141167 116638 141967 6 mem_addr[14]
port 73 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 mem_addr[15]
port 74 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 mem_addr[16]
port 75 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 mem_addr[17]
port 76 nsew signal output
rlabel metal2 s 22558 141167 22614 141967 6 mem_addr[18]
port 77 nsew signal output
rlabel metal3 s 139023 54408 139823 54528 6 mem_addr[19]
port 78 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 mem_addr[1]
port 79 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 mem_addr[20]
port 80 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 mem_addr[21]
port 81 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 mem_addr[22]
port 82 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 mem_addr[23]
port 83 nsew signal output
rlabel metal2 s 76010 141167 76066 141967 6 mem_addr[24]
port 84 nsew signal output
rlabel metal3 s 139023 47608 139823 47728 6 mem_addr[25]
port 85 nsew signal output
rlabel metal3 s 139023 34688 139823 34808 6 mem_addr[26]
port 86 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 mem_addr[27]
port 87 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 mem_addr[28]
port 88 nsew signal output
rlabel metal2 s 36082 141167 36138 141967 6 mem_addr[29]
port 89 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 mem_addr[2]
port 90 nsew signal output
rlabel metal3 s 139023 58488 139823 58608 6 mem_addr[30]
port 91 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 mem_addr[31]
port 92 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 mem_addr[3]
port 93 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 mem_addr[4]
port 94 nsew signal output
rlabel metal2 s 83094 141167 83150 141967 6 mem_addr[5]
port 95 nsew signal output
rlabel metal2 s 7746 141167 7802 141967 6 mem_addr[6]
port 96 nsew signal output
rlabel metal3 s 139023 128528 139823 128648 6 mem_addr[7]
port 97 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 mem_addr[8]
port 98 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 mem_addr[9]
port 99 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 mem_instr
port 100 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 mem_la_addr[0]
port 101 nsew signal output
rlabel metal3 s 139023 76848 139823 76968 6 mem_la_addr[10]
port 102 nsew signal output
rlabel metal2 s 662 141167 718 141967 6 mem_la_addr[11]
port 103 nsew signal output
rlabel metal2 s 47674 141167 47730 141967 6 mem_la_addr[12]
port 104 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 mem_la_addr[13]
port 105 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 mem_la_addr[14]
port 106 nsew signal output
rlabel metal2 s 89534 141167 89590 141967 6 mem_la_addr[15]
port 107 nsew signal output
rlabel metal3 s 139023 97248 139823 97368 6 mem_la_addr[16]
port 108 nsew signal output
rlabel metal2 s 1950 141167 2006 141967 6 mem_la_addr[17]
port 109 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 mem_la_addr[18]
port 110 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 mem_la_addr[19]
port 111 nsew signal output
rlabel metal3 s 139023 24488 139823 24608 6 mem_la_addr[1]
port 112 nsew signal output
rlabel metal2 s 5170 141167 5226 141967 6 mem_la_addr[20]
port 113 nsew signal output
rlabel metal2 s 61198 141167 61254 141967 6 mem_la_addr[21]
port 114 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 mem_la_addr[22]
port 115 nsew signal output
rlabel metal2 s 28998 141167 29054 141967 6 mem_la_addr[23]
port 116 nsew signal output
rlabel metal2 s 19982 141167 20038 141967 6 mem_la_addr[24]
port 117 nsew signal output
rlabel metal3 s 139023 119688 139823 119808 6 mem_la_addr[25]
port 118 nsew signal output
rlabel metal2 s 18694 141167 18750 141967 6 mem_la_addr[26]
port 119 nsew signal output
rlabel metal3 s 139023 30608 139823 30728 6 mem_la_addr[27]
port 120 nsew signal output
rlabel metal2 s 9034 141167 9090 141967 6 mem_la_addr[28]
port 121 nsew signal output
rlabel metal3 s 139023 131248 139823 131368 6 mem_la_addr[29]
port 122 nsew signal output
rlabel metal3 s 139023 51688 139823 51808 6 mem_la_addr[2]
port 123 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 mem_la_addr[30]
port 124 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 mem_la_addr[31]
port 125 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 mem_la_addr[3]
port 126 nsew signal output
rlabel metal3 s 139023 114248 139823 114368 6 mem_la_addr[4]
port 127 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 mem_la_addr[5]
port 128 nsew signal output
rlabel metal3 s 139023 116968 139823 117088 6 mem_la_addr[6]
port 129 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 mem_la_addr[7]
port 130 nsew signal output
rlabel metal3 s 139023 27208 139823 27328 6 mem_la_addr[8]
port 131 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 mem_la_addr[9]
port 132 nsew signal output
rlabel metal3 s 139023 31968 139823 32088 6 mem_la_read
port 133 nsew signal output
rlabel metal2 s 123022 141167 123078 141967 6 mem_la_wdata[0]
port 134 nsew signal output
rlabel metal3 s 139023 101328 139823 101448 6 mem_la_wdata[10]
port 135 nsew signal output
rlabel metal2 s 68282 141167 68338 141967 6 mem_la_wdata[11]
port 136 nsew signal output
rlabel metal2 s 25134 141167 25190 141967 6 mem_la_wdata[12]
port 137 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 mem_la_wdata[13]
port 138 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 mem_la_wdata[14]
port 139 nsew signal output
rlabel metal2 s 54758 141167 54814 141967 6 mem_la_wdata[15]
port 140 nsew signal output
rlabel metal2 s 115294 141167 115350 141967 6 mem_la_wdata[16]
port 141 nsew signal output
rlabel metal2 s 128818 141167 128874 141967 6 mem_la_wdata[17]
port 142 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 mem_la_wdata[18]
port 143 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 mem_la_wdata[19]
port 144 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 mem_la_wdata[1]
port 145 nsew signal output
rlabel metal3 s 139023 99968 139823 100088 6 mem_la_wdata[20]
port 146 nsew signal output
rlabel metal3 s 139023 81608 139823 81728 6 mem_la_wdata[21]
port 147 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 mem_la_wdata[22]
port 148 nsew signal output
rlabel metal3 s 139023 98608 139823 98728 6 mem_la_wdata[23]
port 149 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 mem_la_wdata[24]
port 150 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 mem_la_wdata[25]
port 151 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 mem_la_wdata[26]
port 152 nsew signal output
rlabel metal2 s 95330 141167 95386 141967 6 mem_la_wdata[27]
port 153 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 mem_la_wdata[28]
port 154 nsew signal output
rlabel metal2 s 59910 141167 59966 141967 6 mem_la_wdata[29]
port 155 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 mem_la_wdata[2]
port 156 nsew signal output
rlabel metal3 s 139023 40128 139823 40248 6 mem_la_wdata[30]
port 157 nsew signal output
rlabel metal2 s 10322 141167 10378 141967 6 mem_la_wdata[31]
port 158 nsew signal output
rlabel metal3 s 139023 33328 139823 33448 6 mem_la_wdata[3]
port 159 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 mem_la_wdata[4]
port 160 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 mem_la_wdata[5]
port 161 nsew signal output
rlabel metal3 s 139023 138048 139823 138168 6 mem_la_wdata[6]
port 162 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 mem_la_wdata[7]
port 163 nsew signal output
rlabel metal3 s 139023 123768 139823 123888 6 mem_la_wdata[8]
port 164 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 mem_la_wdata[9]
port 165 nsew signal output
rlabel metal3 s 139023 61888 139823 62008 6 mem_la_write
port 166 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 mem_la_wstrb[0]
port 167 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 mem_la_wstrb[1]
port 168 nsew signal output
rlabel metal2 s 100482 141167 100538 141967 6 mem_la_wstrb[2]
port 169 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 mem_la_wstrb[3]
port 170 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 mem_rdata[0]
port 171 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 mem_rdata[10]
port 172 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 mem_rdata[11]
port 173 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 mem_rdata[12]
port 174 nsew signal input
rlabel metal2 s 31574 141167 31630 141967 6 mem_rdata[13]
port 175 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 mem_rdata[14]
port 176 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 mem_rdata[15]
port 177 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 mem_rdata[16]
port 178 nsew signal input
rlabel metal3 s 139023 53048 139823 53168 6 mem_rdata[17]
port 179 nsew signal input
rlabel metal2 s 26422 141167 26478 141967 6 mem_rdata[18]
port 180 nsew signal input
rlabel metal2 s 72146 141167 72202 141967 6 mem_rdata[19]
port 181 nsew signal input
rlabel metal2 s 73434 141167 73490 141967 6 mem_rdata[1]
port 182 nsew signal input
rlabel metal3 s 139023 111528 139823 111648 6 mem_rdata[20]
port 183 nsew signal input
rlabel metal2 s 57334 141167 57390 141967 6 mem_rdata[21]
port 184 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 mem_rdata[22]
port 185 nsew signal input
rlabel metal2 s 69570 141167 69626 141967 6 mem_rdata[23]
port 186 nsew signal input
rlabel metal2 s 114006 141167 114062 141967 6 mem_rdata[24]
port 187 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 mem_rdata[25]
port 188 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 mem_rdata[26]
port 189 nsew signal input
rlabel metal2 s 104346 141167 104402 141967 6 mem_rdata[27]
port 190 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 mem_rdata[28]
port 191 nsew signal input
rlabel metal2 s 124310 141167 124366 141967 6 mem_rdata[29]
port 192 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 mem_rdata[2]
port 193 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 mem_rdata[30]
port 194 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 mem_rdata[31]
port 195 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 mem_rdata[3]
port 196 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 mem_rdata[4]
port 197 nsew signal input
rlabel metal2 s 52182 141167 52238 141967 6 mem_rdata[5]
port 198 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 mem_rdata[6]
port 199 nsew signal input
rlabel metal3 s 139023 20408 139823 20528 6 mem_rdata[7]
port 200 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 mem_rdata[8]
port 201 nsew signal input
rlabel metal2 s 80518 141167 80574 141967 6 mem_rdata[9]
port 202 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 mem_ready
port 203 nsew signal input
rlabel metal3 s 139023 50328 139823 50448 6 mem_valid
port 204 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 mem_wdata[0]
port 205 nsew signal output
rlabel metal2 s 53470 141167 53526 141967 6 mem_wdata[10]
port 206 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 mem_wdata[11]
port 207 nsew signal output
rlabel metal2 s 15474 141167 15530 141967 6 mem_wdata[12]
port 208 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 mem_wdata[13]
port 209 nsew signal output
rlabel metal3 s 139023 115608 139823 115728 6 mem_wdata[14]
port 210 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 mem_wdata[15]
port 211 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 mem_wdata[16]
port 212 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 mem_wdata[17]
port 213 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 mem_wdata[18]
port 214 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 mem_wdata[19]
port 215 nsew signal output
rlabel metal2 s 88246 141167 88302 141967 6 mem_wdata[1]
port 216 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 mem_wdata[20]
port 217 nsew signal output
rlabel metal2 s 84382 141167 84438 141967 6 mem_wdata[21]
port 218 nsew signal output
rlabel metal3 s 139023 11568 139823 11688 6 mem_wdata[22]
port 219 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 mem_wdata[23]
port 220 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 mem_wdata[24]
port 221 nsew signal output
rlabel metal3 s 0 121728 800 121848 6 mem_wdata[25]
port 222 nsew signal output
rlabel metal3 s 139023 92488 139823 92608 6 mem_wdata[26]
port 223 nsew signal output
rlabel metal2 s 64418 141167 64474 141967 6 mem_wdata[27]
port 224 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 mem_wdata[28]
port 225 nsew signal output
rlabel metal2 s 111430 141167 111486 141967 6 mem_wdata[29]
port 226 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 mem_wdata[2]
port 227 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 mem_wdata[30]
port 228 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 mem_wdata[31]
port 229 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 mem_wdata[3]
port 230 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 mem_wdata[4]
port 231 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 mem_wdata[5]
port 232 nsew signal output
rlabel metal3 s 139023 6128 139823 6248 6 mem_wdata[6]
port 233 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 mem_wdata[7]
port 234 nsew signal output
rlabel metal2 s 137834 141167 137890 141967 6 mem_wdata[8]
port 235 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 mem_wdata[9]
port 236 nsew signal output
rlabel metal3 s 139023 63248 139823 63368 6 mem_wstrb[0]
port 237 nsew signal output
rlabel metal3 s 139023 48968 139823 49088 6 mem_wstrb[1]
port 238 nsew signal output
rlabel metal3 s 139023 95888 139823 96008 6 mem_wstrb[2]
port 239 nsew signal output
rlabel metal3 s 139023 75488 139823 75608 6 mem_wstrb[3]
port 240 nsew signal output
rlabel metal2 s 6458 141167 6514 141967 6 pcpi_insn[0]
port 241 nsew signal output
rlabel metal3 s 139023 78888 139823 79008 6 pcpi_insn[10]
port 242 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 pcpi_insn[11]
port 243 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 pcpi_insn[12]
port 244 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 pcpi_insn[13]
port 245 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 pcpi_insn[14]
port 246 nsew signal output
rlabel metal2 s 14186 141167 14242 141967 6 pcpi_insn[15]
port 247 nsew signal output
rlabel metal3 s 139023 7488 139823 7608 6 pcpi_insn[16]
port 248 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 pcpi_insn[17]
port 249 nsew signal output
rlabel metal2 s 132682 141167 132738 141967 6 pcpi_insn[18]
port 250 nsew signal output
rlabel metal2 s 62486 141167 62542 141967 6 pcpi_insn[19]
port 251 nsew signal output
rlabel metal2 s 108210 141167 108266 141967 6 pcpi_insn[1]
port 252 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 pcpi_insn[20]
port 253 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 pcpi_insn[21]
port 254 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 pcpi_insn[22]
port 255 nsew signal output
rlabel metal2 s 99194 141167 99250 141967 6 pcpi_insn[23]
port 256 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 pcpi_insn[24]
port 257 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 pcpi_insn[25]
port 258 nsew signal output
rlabel metal3 s 139023 132608 139823 132728 6 pcpi_insn[26]
port 259 nsew signal output
rlabel metal3 s 139023 139408 139823 139528 6 pcpi_insn[27]
port 260 nsew signal output
rlabel metal3 s 139023 118328 139823 118448 6 pcpi_insn[28]
port 261 nsew signal output
rlabel metal2 s 65706 141167 65762 141967 6 pcpi_insn[29]
port 262 nsew signal output
rlabel metal3 s 139023 112888 139823 113008 6 pcpi_insn[2]
port 263 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 pcpi_insn[30]
port 264 nsew signal output
rlabel metal2 s 127530 141167 127586 141967 6 pcpi_insn[31]
port 265 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 pcpi_insn[3]
port 266 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 pcpi_insn[4]
port 267 nsew signal output
rlabel metal2 s 23846 141167 23902 141967 6 pcpi_insn[5]
port 268 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 pcpi_insn[6]
port 269 nsew signal output
rlabel metal3 s 139023 688 139823 808 6 pcpi_insn[7]
port 270 nsew signal output
rlabel metal2 s 136546 141167 136602 141967 6 pcpi_insn[8]
port 271 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 pcpi_insn[9]
port 272 nsew signal output
rlabel metal2 s 56046 141167 56102 141967 6 pcpi_rd[0]
port 273 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 pcpi_rd[10]
port 274 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 pcpi_rd[11]
port 275 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 pcpi_rd[12]
port 276 nsew signal input
rlabel metal2 s 119158 141167 119214 141967 6 pcpi_rd[13]
port 277 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 pcpi_rd[14]
port 278 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 pcpi_rd[15]
port 279 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 pcpi_rd[16]
port 280 nsew signal input
rlabel metal3 s 139023 65968 139823 66088 6 pcpi_rd[17]
port 281 nsew signal input
rlabel metal3 s 139023 91128 139823 91248 6 pcpi_rd[18]
port 282 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 pcpi_rd[19]
port 283 nsew signal input
rlabel metal2 s 49606 141167 49662 141967 6 pcpi_rd[1]
port 284 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 pcpi_rd[20]
port 285 nsew signal input
rlabel metal3 s 139023 87048 139823 87168 6 pcpi_rd[21]
port 286 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 pcpi_rd[22]
port 287 nsew signal input
rlabel metal3 s 139023 70048 139823 70168 6 pcpi_rd[23]
port 288 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 pcpi_rd[24]
port 289 nsew signal input
rlabel metal2 s 126242 141167 126298 141967 6 pcpi_rd[25]
port 290 nsew signal input
rlabel metal3 s 139023 10208 139823 10328 6 pcpi_rd[26]
port 291 nsew signal input
rlabel metal2 s 86958 141167 87014 141967 6 pcpi_rd[27]
port 292 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 pcpi_rd[28]
port 293 nsew signal input
rlabel metal2 s 38658 141167 38714 141967 6 pcpi_rd[29]
port 294 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 pcpi_rd[2]
port 295 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 pcpi_rd[30]
port 296 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 pcpi_rd[31]
port 297 nsew signal input
rlabel metal3 s 139023 89768 139823 89888 6 pcpi_rd[3]
port 298 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 pcpi_rd[4]
port 299 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 pcpi_rd[5]
port 300 nsew signal input
rlabel metal2 s 45098 141167 45154 141967 6 pcpi_rd[6]
port 301 nsew signal input
rlabel metal2 s 121734 141167 121790 141967 6 pcpi_rd[7]
port 302 nsew signal input
rlabel metal3 s 139023 105408 139823 105528 6 pcpi_rd[8]
port 303 nsew signal input
rlabel metal2 s 39946 141167 40002 141967 6 pcpi_rd[9]
port 304 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 pcpi_ready
port 305 nsew signal input
rlabel metal3 s 139023 21768 139823 21888 6 pcpi_rs1[0]
port 306 nsew signal output
rlabel metal2 s 30286 141167 30342 141967 6 pcpi_rs1[10]
port 307 nsew signal output
rlabel metal3 s 139023 46248 139823 46368 6 pcpi_rs1[11]
port 308 nsew signal output
rlabel metal2 s 96618 141167 96674 141967 6 pcpi_rs1[12]
port 309 nsew signal output
rlabel metal2 s 66994 141167 67050 141967 6 pcpi_rs1[13]
port 310 nsew signal output
rlabel metal2 s 12898 141167 12954 141967 6 pcpi_rs1[14]
port 311 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 pcpi_rs1[15]
port 312 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 pcpi_rs1[16]
port 313 nsew signal output
rlabel metal3 s 139023 102688 139823 102808 6 pcpi_rs1[17]
port 314 nsew signal output
rlabel metal3 s 139023 94528 139823 94648 6 pcpi_rs1[18]
port 315 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 pcpi_rs1[19]
port 316 nsew signal output
rlabel metal3 s 139023 82968 139823 83088 6 pcpi_rs1[1]
port 317 nsew signal output
rlabel metal3 s 139023 41488 139823 41608 6 pcpi_rs1[20]
port 318 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 pcpi_rs1[21]
port 319 nsew signal output
rlabel metal2 s 92110 141167 92166 141967 6 pcpi_rs1[22]
port 320 nsew signal output
rlabel metal2 s 131394 141167 131450 141967 6 pcpi_rs1[23]
port 321 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 pcpi_rs1[24]
port 322 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 pcpi_rs1[25]
port 323 nsew signal output
rlabel metal3 s 139023 29248 139823 29368 6 pcpi_rs1[26]
port 324 nsew signal output
rlabel metal2 s 21270 141167 21326 141967 6 pcpi_rs1[27]
port 325 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 pcpi_rs1[28]
port 326 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 pcpi_rs1[29]
port 327 nsew signal output
rlabel metal2 s 50894 141167 50950 141967 6 pcpi_rs1[2]
port 328 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 pcpi_rs1[30]
port 329 nsew signal output
rlabel metal3 s 139023 135328 139823 135448 6 pcpi_rs1[31]
port 330 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 pcpi_rs1[3]
port 331 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 pcpi_rs1[4]
port 332 nsew signal output
rlabel metal3 s 139023 57128 139823 57248 6 pcpi_rs1[5]
port 333 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 pcpi_rs1[6]
port 334 nsew signal output
rlabel metal2 s 110142 141167 110198 141967 6 pcpi_rs1[7]
port 335 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 pcpi_rs1[8]
port 336 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 pcpi_rs1[9]
port 337 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 pcpi_rs2[0]
port 338 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 pcpi_rs2[10]
port 339 nsew signal output
rlabel metal3 s 139023 36048 139823 36168 6 pcpi_rs2[11]
port 340 nsew signal output
rlabel metal2 s 46386 141167 46442 141967 6 pcpi_rs2[12]
port 341 nsew signal output
rlabel metal3 s 139023 122408 139823 122528 6 pcpi_rs2[13]
port 342 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 pcpi_rs2[14]
port 343 nsew signal output
rlabel metal3 s 0 123088 800 123208 6 pcpi_rs2[15]
port 344 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 pcpi_rs2[16]
port 345 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 pcpi_rs2[17]
port 346 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 pcpi_rs2[18]
port 347 nsew signal output
rlabel metal3 s 139023 71408 139823 71528 6 pcpi_rs2[19]
port 348 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 pcpi_rs2[1]
port 349 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 pcpi_rs2[20]
port 350 nsew signal output
rlabel metal2 s 130106 141167 130162 141967 6 pcpi_rs2[21]
port 351 nsew signal output
rlabel metal2 s 11610 141167 11666 141967 6 pcpi_rs2[22]
port 352 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 pcpi_rs2[23]
port 353 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 pcpi_rs2[24]
port 354 nsew signal output
rlabel metal2 s 133970 141167 134026 141967 6 pcpi_rs2[25]
port 355 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 pcpi_rs2[26]
port 356 nsew signal output
rlabel metal3 s 139023 110168 139823 110288 6 pcpi_rs2[27]
port 357 nsew signal output
rlabel metal3 s 139023 44208 139823 44328 6 pcpi_rs2[28]
port 358 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 pcpi_rs2[29]
port 359 nsew signal output
rlabel metal2 s 117870 141167 117926 141967 6 pcpi_rs2[2]
port 360 nsew signal output
rlabel metal2 s 37370 141167 37426 141967 6 pcpi_rs2[30]
port 361 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 pcpi_rs2[31]
port 362 nsew signal output
rlabel metal3 s 139023 84328 139823 84448 6 pcpi_rs2[3]
port 363 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 pcpi_rs2[4]
port 364 nsew signal output
rlabel metal3 s 139023 38768 139823 38888 6 pcpi_rs2[5]
port 365 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 pcpi_rs2[6]
port 366 nsew signal output
rlabel metal3 s 139023 2048 139823 2168 6 pcpi_rs2[7]
port 367 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 pcpi_rs2[8]
port 368 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 pcpi_rs2[9]
port 369 nsew signal output
rlabel metal3 s 139023 59848 139823 59968 6 pcpi_valid
port 370 nsew signal output
rlabel metal2 s 112718 141167 112774 141967 6 pcpi_wait
port 371 nsew signal input
rlabel metal3 s 139023 127168 139823 127288 6 pcpi_wr
port 372 nsew signal input
rlabel metal3 s 139023 4768 139823 4888 6 resetn
port 373 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 trace_data[0]
port 374 nsew signal output
rlabel metal3 s 139023 80248 139823 80368 6 trace_data[10]
port 375 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 trace_data[11]
port 376 nsew signal output
rlabel metal3 s 139023 129888 139823 130008 6 trace_data[12]
port 377 nsew signal output
rlabel metal2 s 106922 141167 106978 141967 6 trace_data[13]
port 378 nsew signal output
rlabel metal3 s 139023 13608 139823 13728 6 trace_data[14]
port 379 nsew signal output
rlabel metal2 s 101770 141167 101826 141967 6 trace_data[15]
port 380 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 trace_data[16]
port 381 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 trace_data[17]
port 382 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 trace_data[18]
port 383 nsew signal output
rlabel metal2 s 18 0 74 800 6 trace_data[19]
port 384 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 trace_data[1]
port 385 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 trace_data[20]
port 386 nsew signal output
rlabel metal3 s 0 125808 800 125928 6 trace_data[21]
port 387 nsew signal output
rlabel metal2 s 41234 141167 41290 141967 6 trace_data[22]
port 388 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 trace_data[23]
port 389 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 trace_data[24]
port 390 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 trace_data[25]
port 391 nsew signal output
rlabel metal2 s 74722 141167 74778 141967 6 trace_data[26]
port 392 nsew signal output
rlabel metal2 s 43810 141167 43866 141967 6 trace_data[27]
port 393 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 trace_data[28]
port 394 nsew signal output
rlabel metal2 s 97906 141167 97962 141967 6 trace_data[29]
port 395 nsew signal output
rlabel metal3 s 139023 37408 139823 37528 6 trace_data[2]
port 396 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 trace_data[30]
port 397 nsew signal output
rlabel metal3 s 139023 108128 139823 108248 6 trace_data[31]
port 398 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 trace_data[32]
port 399 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 trace_data[33]
port 400 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 trace_data[34]
port 401 nsew signal output
rlabel metal3 s 139023 104048 139823 104168 6 trace_data[35]
port 402 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 trace_data[3]
port 403 nsew signal output
rlabel metal2 s 93398 141167 93454 141967 6 trace_data[4]
port 404 nsew signal output
rlabel metal2 s 90822 141167 90878 141967 6 trace_data[5]
port 405 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 trace_data[6]
port 406 nsew signal output
rlabel metal2 s 16762 141167 16818 141967 6 trace_data[7]
port 407 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 trace_data[8]
port 408 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 trace_data[9]
port 409 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 trace_valid
port 410 nsew signal output
rlabel metal3 s 139023 68688 139823 68808 6 trap
port 411 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 139823 141967
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 55707800
string GDS_FILE /home/aanujdu/z2a/caravel_user_project/openlane/picorv32a/runs/picorv32a/results/finishing/picorv32a.magic.gds
string GDS_START 1547148
<< end >>

